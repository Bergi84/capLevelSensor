-- megafunction wizard: %ALTIOBUF%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: altiobuf_bidir 

-- ============================================================
-- File Name: ioBuf.vhd
-- Megafunction Name(s):
-- 			altiobuf_bidir
--
-- Simulation Library Files(s):
-- 			cycloneive
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 21.1.0 Build 842 10/21/2021 SJ Lite Edition
-- ************************************************************


--Copyright (C) 2021  Intel Corporation. All rights reserved.
--Your use of Intel Corporation's design tools, logic functions 
--and other software and tools, and any partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Intel Program License 
--Subscription Agreement, the Intel Quartus Prime License Agreement,
--the Intel FPGA IP License Agreement, or other applicable license
--agreement, including, without limitation, that your use is for
--the sole purpose of programming logic devices manufactured by
--Intel and sold by Intel or its authorized distributors.  Please
--refer to the applicable agreement for further details, at
--https://fpgasoftware.intel.com/eula.


--altiobuf_bidir CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone IV E" ENABLE_BUS_HOLD="FALSE" NUMBER_OF_CHANNELS=4 OPEN_DRAIN_OUTPUT="FALSE" USE_DIFFERENTIAL_MODE="FALSE" USE_DYNAMIC_TERMINATION_CONTROL="FALSE" USE_TERMINATION_CONTROL="FALSE" datain dataio dataout oe
--VERSION_BEGIN 21.1 cbx_altiobuf_bidir 2021:10:21:11:03:22:SJ cbx_mgl 2021:10:21:11:03:46:SJ cbx_stratixiii 2021:10:21:11:03:22:SJ cbx_stratixv 2021:10:21:11:03:22:SJ  VERSION_END

 LIBRARY cycloneive;
 USE cycloneive.all;

--synthesis_resources = cycloneive_io_ibuf 4 cycloneive_io_obuf 4 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  ioBuf_iobuf_bidir_60p IS 
	 PORT 
	 ( 
		 datain	:	IN  STD_LOGIC_VECTOR (3 DOWNTO 0);
		 dataio	:	INOUT  STD_LOGIC_VECTOR (3 DOWNTO 0);
		 dataout	:	OUT  STD_LOGIC_VECTOR (3 DOWNTO 0);
		 oe	:	IN  STD_LOGIC_VECTOR (3 DOWNTO 0)
	 ); 
 END ioBuf_iobuf_bidir_60p;

 ARCHITECTURE RTL OF ioBuf_iobuf_bidir_60p IS

	 SIGNAL  wire_ibufa_i	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_ibufa_o	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_obufa_i	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_obufa_o	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_obufa_oe	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 COMPONENT  cycloneive_io_ibuf
	 GENERIC 
	 (
		bus_hold	:	STRING := "false";
		differential_mode	:	STRING := "false";
		simulate_z_as	:	STRING := "Z";
		lpm_type	:	STRING := "cycloneive_io_ibuf"
	 );
	 PORT
	 ( 
		i	:	IN STD_LOGIC := '0';
		ibar	:	IN STD_LOGIC := '0';
		o	:	OUT STD_LOGIC
	 ); 
	 END COMPONENT;
	 COMPONENT  cycloneive_io_obuf
	 GENERIC 
	 (
		bus_hold	:	STRING := "false";
		open_drain_output	:	STRING := "false";
		lpm_type	:	STRING := "cycloneive_io_obuf"
	 );
	 PORT
	 ( 
		i	:	IN STD_LOGIC := '0';
		o	:	OUT STD_LOGIC;
		obar	:	OUT STD_LOGIC;
		oe	:	IN STD_LOGIC := '1';
		seriesterminationcontrol	:	IN STD_LOGIC_VECTOR(15 DOWNTO 0) := (OTHERS => '0')
	 ); 
	 END COMPONENT;
 BEGIN

	dataio <= wire_obufa_o;
	dataout <= wire_ibufa_o;
	wire_ibufa_i <= dataio;
	loop0 : FOR i IN 0 TO 3 GENERATE 
	  ibufa :  cycloneive_io_ibuf
	  GENERIC MAP (
		bus_hold => "false",
		differential_mode => "false"
	  )
	  PORT MAP ( 
		i => wire_ibufa_i(i),
		o => wire_ibufa_o(i)
	  );
	END GENERATE loop0;
	wire_obufa_i <= datain;
	wire_obufa_oe <= oe;
	loop1 : FOR i IN 0 TO 3 GENERATE 
	  obufa :  cycloneive_io_obuf
	  GENERIC MAP (
		bus_hold => "false",
		open_drain_output => "false"
	  )
	  PORT MAP ( 
		i => wire_obufa_i(i),
		o => wire_obufa_o(i),
		oe => wire_obufa_oe(i)
	  );
	END GENERATE loop1;

 END RTL; --ioBuf_iobuf_bidir_60p
--VALID FILE


LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY ioBuf IS
	PORT
	(
		datain		: IN STD_LOGIC_VECTOR (3 DOWNTO 0);
		oe		: IN STD_LOGIC_VECTOR (3 DOWNTO 0);
		dataio		: INOUT STD_LOGIC_VECTOR (3 DOWNTO 0);
		dataout		: OUT STD_LOGIC_VECTOR (3 DOWNTO 0)
	);
END ioBuf;


ARCHITECTURE RTL OF iobuf IS

	SIGNAL sub_wire0	: STD_LOGIC_VECTOR (3 DOWNTO 0);



	COMPONENT ioBuf_iobuf_bidir_60p
	PORT (
			datain	: IN STD_LOGIC_VECTOR (3 DOWNTO 0);
			oe	: IN STD_LOGIC_VECTOR (3 DOWNTO 0);
			dataout	: OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
			dataio	: INOUT STD_LOGIC_VECTOR (3 DOWNTO 0)
	);
	END COMPONENT;

BEGIN
	dataout    <= sub_wire0(3 DOWNTO 0);

	ioBuf_iobuf_bidir_60p_component : ioBuf_iobuf_bidir_60p
	PORT MAP (
		datain => datain,
		oe => oe,
		dataout => sub_wire0,
		dataio => dataio
	);



END RTL;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone IV E"
-- Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
-- Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
-- Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Cyclone IV E"
-- Retrieval info: CONSTANT: enable_bus_hold STRING "FALSE"
-- Retrieval info: CONSTANT: number_of_channels NUMERIC "4"
-- Retrieval info: CONSTANT: open_drain_output STRING "FALSE"
-- Retrieval info: CONSTANT: use_differential_mode STRING "FALSE"
-- Retrieval info: CONSTANT: use_dynamic_termination_control STRING "FALSE"
-- Retrieval info: CONSTANT: use_termination_control STRING "FALSE"
-- Retrieval info: USED_PORT: datain 0 0 4 0 INPUT NODEFVAL "datain[3..0]"
-- Retrieval info: USED_PORT: dataio 0 0 4 0 BIDIR NODEFVAL "dataio[3..0]"
-- Retrieval info: USED_PORT: dataout 0 0 4 0 OUTPUT NODEFVAL "dataout[3..0]"
-- Retrieval info: USED_PORT: oe 0 0 4 0 INPUT NODEFVAL "oe[3..0]"
-- Retrieval info: CONNECT: @datain 0 0 4 0 datain 0 0 4 0
-- Retrieval info: CONNECT: @oe 0 0 4 0 oe 0 0 4 0
-- Retrieval info: CONNECT: dataio 0 0 4 0 @dataio 0 0 4 0
-- Retrieval info: CONNECT: dataout 0 0 4 0 @dataout 0 0 4 0
-- Retrieval info: GEN_FILE: TYPE_NORMAL ioBuf.vhd TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL ioBuf.inc FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL ioBuf.cmp TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL ioBuf.bsf FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL ioBuf_inst.vhd FALSE
-- Retrieval info: LIB_FILE: cycloneive
